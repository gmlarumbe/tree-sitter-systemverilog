module a ();

always @(posedge clk, negedge rst_n) begin end

endmodule
