`some_macro(arg1)
