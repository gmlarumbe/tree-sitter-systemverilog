  parameter int AW = -1;
