// Section 140.2: $fopen and $fclose

fd = $fopen ("file_name", "rb+"); // open for update (reading and writing)


