initial begin
    cast_t1 temp1;
    cast_t2 temp2;
    temp1 = expr_1;
    temp2 = expr_2;
    A = temp1 + temp2;
end
