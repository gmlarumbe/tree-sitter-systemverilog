module mod ();
  always_comb foo = bar.baz.bat[7:0];
endmodule
