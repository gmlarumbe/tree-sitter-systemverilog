// Section 120.1: `timescale
 
`timescale 10ns / 1ps


