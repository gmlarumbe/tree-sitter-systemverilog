// Section 106.3: Typedef

typedef union { int X; shortreal Y; } FloatingPoint; 
FloatingPoint N;
N.Y = 0.0; 


