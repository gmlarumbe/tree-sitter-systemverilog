// Section 8.6: Attribute

// Attribute attached to a module definition
(* optimize_power *) module M1 (/*...*/); endmodule


