module mod ();
  assign a = b[1];
endmodule
