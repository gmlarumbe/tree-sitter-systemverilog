task foo(input logic in, output logic out);
     foo = foo2;
endtask
