// Section 2.4: Always
  
always_latch
  if (Enable) Q <= D;


