module test;
    initial $monitor("%d, %d, %d", a, b, c);
endmodule
