function void foo;
    a = package_scope::class_type::member[a].a().method();
endfunction
