function void foo();
    a = this.a.b.c(.arg1(arg1), .arg2(arg2));
endfunction
