function void foo();
    this.in_use[i+1].get_start_offset();
endfunction
