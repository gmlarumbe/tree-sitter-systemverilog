function void foo();
    a = init();
endfunction
