module mod;
endmodule
