module mod #(
  parameter A=5,
  parameter B=10
)();

endmodule
