class foo;

    extern function void foo;
    extern task  foo2;

endclass
