EMPTY <= #`TCQ 1'b1;
