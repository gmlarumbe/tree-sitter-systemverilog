module x;
    always begin
        a <= {5{1'b0}};
    end
endmodule
