// hierarchical identifier with constant expressions plus select
function f;
    left.member[0].nested[1] = right.member[0].nested[1];
endfunction
