function void class_scope::method(some_type arg);
    foo = foo2;
endfunction : method
