class class_name;
  data members;  // class properties

  // class methods
  function function_name;
  // . . .
  endfunction

  task task_name;
  // . . .
  endtask
endclass
