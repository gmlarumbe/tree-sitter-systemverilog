// Section 40.1: Force

initial begin
    force f = a && b;
    /*...*/
    release f;
end


