// Section 142.1: $monitor

initial
  $monitor("%t : a = %b, f = %b", $realtime, a, f);


