function void foo;
  `MY_MACRO.method_call();
endfunction
