`undefineall
