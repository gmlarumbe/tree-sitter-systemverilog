module mod #(
  parameter type T=logic,
  parameter type Q=bit
)();

endmodule
