function void foo();
    if (callbacks.size()) begin
        return;
    end
endfunction
