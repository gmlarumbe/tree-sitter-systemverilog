// Section 76.4: Parameter

// Named association of parameters
module UseShifter(/*...*/);
  Shifter #(.Nbits(10)) MyDecadeShifter(/*...*/);
endmodule


