`define_var


