module foo;

    logic       data0 [*];
    logic       data1 [int];
    logic       data2 [string];
    logic [3:0] data3 [logic];
    int         data3 [bit[3:0]];

endmodule;
