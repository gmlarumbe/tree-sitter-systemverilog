// hierarchical identifier with non-constant expressions (i++) plus select
function f;
    left.member[i++].nested[1] = right.member[i++].nested[1];
endfunction
