function f;
    left.member[1][2] = right.member[1][2];
endfunction
