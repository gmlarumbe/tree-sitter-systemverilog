module mod ();
  always_comb foo = bar.baz[7:0];
endmodule
