a.a.a = a.a.a[a] + a.a.a[a];
a.a.a = (a.a.a[a] + a.a.a[a]);
a.a.a = ~(a.a.a[a] + a.a.a[a]);
a.a.a = a.a.a[0] + a.a.a[0];
a.a.a = (a.a.a[0] + a.a.a[0]);
a.a.a = ~(a.a.a[0] + a.a.a[0]);
a.a.a = a.a.a[a+0] + a.a.a[a+0] ;
a.a.a = (a.a.a[a+0] + a.a.a[a+0]) ;
a.a.a = ~(a.a.a[a+0] + a.a.a[a+0]) ;
a.a.a = a.a.a[0+1] + a.a.a[0+1] ;
a.a.a = (a.a.a[0+1] + a.a.a[0+1]) ;
a.a.a = ~(a.a.a[0+1] + a.a.a[0+1]) ;

a.a.a = a.a.a[a] + a.a.a[a] + a.a.a[a];
a.a.a = (a.a.a[a] + a.a.a[a] + a.a.a[a]);
a.a.a = ~(a.a.a[a] + a.a.a[a] + a.a.a[a]);
a.a.a = a.a.a[0] + a.a.a[0] + a.a.a[0];
a.a.a = (a.a.a[0] + a.a.a[0] + a.a.a[0]);
a.a.a = ~(a.a.a[0] + a.a.a[0] + a.a.a[0]);
a.a.a = a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0];
a.a.a = (a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0]);
a.a.a = ~(a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0]);
a.a.a = a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1];
a.a.a = (a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1]);
a.a.a = ~(a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1]);

a.a.a = a.a.a[a] + a.a.a[a] + a.a.a[a] + a.a.a[a];
a.a.a = (a.a.a[a] + a.a.a[a] + a.a.a[a] + a.a.a[a]);
a.a.a = ~(a.a.a[a] + a.a.a[a] + a.a.a[a] + a.a.a[a]);
a.a.a = a.a.a[0] + a.a.a[0] + a.a.a[0] + a.a.a[a];
a.a.a = (a.a.a[0] + a.a.a[0] + a.a.a[0] + a.a.a[0]);
a.a.a = ~(a.a.a[0] + a.a.a[0] + a.a.a[0] + a.a.a[0]);
a.a.a = a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0];
a.a.a = (a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0]);
a.a.a = ~(a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0] + a.a.a[a+0]);
a.a.a = a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1];
a.a.a = (a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1]);
a.a.a = ~(a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1] + a.a.a[0+1]);
