module mod ();
  wire a;
endmodule
