module mod (output out);
endmodule
