// Section 86.1: Rand

// Random variables in classes
class C;
  rand bit a, b;
endclass

C c = new;

c.randomize();


