bind cpu fpu_props fpu_rules_1(a,b,c);
