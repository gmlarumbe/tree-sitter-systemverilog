// Section 146.1: $timeformat

$timeformat(-10, 2, " x100ps", 20);  // 20.12 x100ps


