// Section 114.1: Wait

wait (count == 10) $display("Count is ten");


