import "DPI-C" context function int foo(string bar);
