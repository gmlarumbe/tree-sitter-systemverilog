function void foo();
    result = this.a.b.c.d.e.f.g.h.i.j.k.l.m.n.o.p.q.r.s.t.u.v.w.x.y.z(.a(1), .b(N-1));
endfunction
