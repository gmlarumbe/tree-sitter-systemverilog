`uvm_do_with(arg, { x == 1; y == 2; });
