module mod ();
  wire a, b, c;
  wire ddd;
  reg ee;
  logic [3:0] fff;
  my_type_t t1, t2;
endmodule
