function void foo();
    init;
endfunction
