package foo;
endpackage
