// Section 131.1: Intersect

// Intersect is used to "and" two sequences, implying a third sequence
assert property (
  a ##1 b ##1 c intersect 1'b1 ##1 d ##1 1'b1 |=> e );


