include *.v;
include ./\*.vg;
