module foo ();

always @(posedge 1'd0) begin end

endmodule
