function void foo;
  `some_macro(arg1)
endfunction
