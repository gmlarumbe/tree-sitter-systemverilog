module mod ();
  assign a = '0;
endmodule
