module abc ();

always_comb
if (foo)
  bar = baz;

endmodule
