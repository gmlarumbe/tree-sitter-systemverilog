// Section 121.1: And (Sequence Operator)

assert property (sig1 and (sig2 ##1 sig3) |-> sig4);


