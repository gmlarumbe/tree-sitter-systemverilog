module x;
    always begin
        lhs <= {(a - b), 1'b0};
    end
endmodule
