module mod #(
  parameter A=5
)();

endmodule
