module abc ();

always begin end
always_ff begin end
always_comb begin end
always_latch begin end

endmodule
