function void foo;
    package_scope::class_type1::class_type2::member[a].a().method();
endfunction
