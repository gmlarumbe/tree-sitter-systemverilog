program foo;
endprogram
