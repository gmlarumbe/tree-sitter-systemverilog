`include "foo.txt"
