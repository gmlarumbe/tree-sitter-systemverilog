module foo;
    logic b;
    assign b = (a.a.a[0] && a.a.a[1]);
endmodule
