module foo;
    specify
        specparam PATHPULSE$clk$q = (0.5,1),
                  PATHPULSE$ = (0.5);
    endspecify
endmodule
