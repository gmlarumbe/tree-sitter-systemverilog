function void foo();
    a = this.fun();
endfunction
