// Section 55.1: Instantiation

// UDP instance
Nand2 (weak1,pull0) #(3,4) (F, A, B);


