initial begin
    if (this.in_use[i] == region) begin
    end
end
