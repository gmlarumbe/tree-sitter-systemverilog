module a_l ();

always begin end

endmodule
