// Section 8.3: Attribute

// Attribute attached to a function call
initial begin
A = add (* mode = "cla" *) (B, C);
end


