// Section 15.4: Class

// Derived class
class ShiftRegister extends Register;
  extern task shiftleft();
  extern task shiftright();
endclass


