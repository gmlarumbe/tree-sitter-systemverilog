module foo;
  block u_block_1 (if1.signal);
  block u_block_2 (if1.signal, if2.signal);
endmodule : foo
