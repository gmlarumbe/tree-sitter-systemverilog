function int foo(string bar, type1 baz);
endfunction
