function f;
    left[i+1][1:0] = right[i+1][1:0];
endfunction
