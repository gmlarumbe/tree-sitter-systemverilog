// Section 54.5: Inside

initial begin
string I;
a = I inside {["abc":"def"]};       // I between "abc" and "def"
end

