bind cpu: cpu1, cpu2, cpu3 fpu_props fpu_rules_1(a, b, c);
