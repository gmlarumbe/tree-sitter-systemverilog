module mod (
  input foo,
  input [3:0] bar,
  output logic [3:0] qux,
  input br_pkt_t dec_i0_brp,
  input wire ham
);

endmodule
