module mod ();
  assign {a, b} = foo;
endmodule
