function void foo();
    a = this.super.fun();
endfunction
