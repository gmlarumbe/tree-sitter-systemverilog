// Section 68.4: Module

// Nested modules
module Mod2(/*...*/);
  module and2(input I1, I2, output O);
    /*...*/
  endmodule
  /*...*/
  and2 U1(/*...*/), U2(/*...*/), U3(/*...*/);
  /*...*/
endmodule


