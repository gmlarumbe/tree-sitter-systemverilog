module mod #(
  parameter  A = 5,
  localparam B = 32/4
)();

endmodule
