module mod ();
  assign a = b;
endmodule
