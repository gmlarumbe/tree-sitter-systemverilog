module mod (clk);
  input clk;
endmodule
