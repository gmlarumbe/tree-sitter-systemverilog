// Section 76.2: Parameter

// Sized parameters
parameter [2:0] Idle = 3'b100, Go1 = 3'b010, Go2 = 3'b001;


