uvm_resource_db#(virtual input_if)::set("env", "input_if", in);
