function f;
    left.member.nested = right.member.nested;
endfunction
