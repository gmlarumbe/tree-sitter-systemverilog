function void foo;
  `MY_MACRO.identifier = 0;
endfunction
