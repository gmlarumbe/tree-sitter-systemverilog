// Section 119.1: `pragma

`pragma resetall
`pragma protect encoding=(enctype="uuencode")
 

