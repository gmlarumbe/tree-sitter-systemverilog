module mod ();
  wire [31:0] a;
endmodule
