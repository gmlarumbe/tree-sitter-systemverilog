`foo(module)
