module mod #(
  parameter type T=logic
)();

endmodule
