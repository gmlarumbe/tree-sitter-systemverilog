// hierarchical identifier with constant expressions plus select and part_select
function f;
    left.member[0].nested[1][2][1:0] = right.member[0].nested[1][2][1:0];
endfunction
