// Section 68.3: Module

module MinMax #(parameter P) (
  input MinMax1,              // ANSI-style port declaration
  input [3:0] X, Y,
  output logic [3:0] Z);
  /*...*/
endmodule


