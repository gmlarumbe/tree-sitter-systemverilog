class comp extends uvm_component;
  `uvm_component_utils(comp)
  // ...
endclass
