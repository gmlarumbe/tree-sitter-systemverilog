`undef Dff
