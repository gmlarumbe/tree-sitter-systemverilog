typedef my_class#(param) my_type_t;
