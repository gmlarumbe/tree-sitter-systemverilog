function void foo;
    class_type::method();
endfunction
