function void foo;
  top.`MY_MACRO.member = 0;
endfunction
