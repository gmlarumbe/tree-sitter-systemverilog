module a ();

always @(posedge clk or negedge rst_n or signal) begin end

endmodule
