`Dff(5, 7)
