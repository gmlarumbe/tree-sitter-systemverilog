function f;
    left.member[1][2][1:0] = right.member[1][2][1:0];
endfunction
