// Section 134.1: Restrict

r1: restrict property (@(posedge clk) mode == 2'b00);


