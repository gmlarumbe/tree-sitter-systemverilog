typedef logic[7:0] byte_t;
