// Section 98.1: String Literal

logic [23:0] MonthName[1:12];

initial
begin
  MonthName[1] =  "Jan";
  MonthName[2]  = "Feb";
  MonthName[3]  = "Mar";
  MonthName[4]  = "Apr";
  MonthName[5]  = "May";
  MonthName[6]  = "Jun";
  MonthName[7]  = "Jul";
  MonthName[8]  = "Aug";
  MonthName[9]  = "Sep";
  MonthName[10] = "Oct";
  MonthName[11] = "Nov";
  MonthName[12] = "Dec";
end


