// Section 38.1: Final

final begin
  $display("Simulation ended: %0d errors.", error_count);
end


