function f;
    left[1][2][1:0] = right[1][3][1:0];
endfunction
