// Section 1.2: Alias

// C is implicitly declared as an 1-bit wire
wire [8:0] word9;
wire [7:0] word;
alias word9 = {word, C};


