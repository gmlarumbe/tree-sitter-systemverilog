typedef package_scope::element my_type_t;
typedef class_type#(param)::element my_type_t;
