module a ();

always @(comb1 or comb2 or comb3 or comb4) begin end

endmodule
