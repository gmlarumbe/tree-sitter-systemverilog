module mod ();
  assign a = b[Param+1:0];
endmodule
