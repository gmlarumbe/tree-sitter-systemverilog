// Section 62.3: Library

// All *.v in this directory and in ../archives belong to library MyDesign
// (uncomment the following to use)
// library MyDesign
//   ./*.v,  // equivalently *.v,
//   ../archives/*.v ;


