// Section 93.1: Statement

LabelA: Statement;
LabelB: begin
  /*...*/
end


