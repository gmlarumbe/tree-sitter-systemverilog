package my_pkg;
    `include "some_file.svh"
endpackage
