// Section 69.2: Name

// Illegal names
logic 123a;                   // Starts with a number
logic $data;                  // Starts with a dollar
logic module;                 // A keyword


