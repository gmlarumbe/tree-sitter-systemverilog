module foo;

    logic       data1 [0:CHANNELS-1];
    logic       data2 [CHANNELS];
    logic [3:0] data3 [CHANNELS];

endmodule;
