// Section 103.1: This

class AClass;
  int Var1;               // Var1 is a property of AClass
  function new (int Var1); // Var1 is an argument of the constructor
    this.Var1 = Var1;     // The instance property is accessed using this
  endfunction
endclass


