function void foo;
   pred = new [predecessors.size()];
endfunction
