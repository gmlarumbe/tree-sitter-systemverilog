virtual class foo;

    virtual function void foo;
    endfunction

endclass
