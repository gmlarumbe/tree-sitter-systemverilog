// Section 101.4: Task

// Argument of type array
task ATask(input [15:0][7:0] A, B[15:0],
           output [15:0][7:0] C[1:0]);
  /*...*/
endtask


