module mod #(
  parameter type T=logic,
                 Q=bit,
  parameter type A = int,
  localparam type D = int
)();

endmodule
