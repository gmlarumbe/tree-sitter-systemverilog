// Section 14.1: Chandle

// Standard C functions imported in SystemVerilog:
import "DPI-C" function chandle malloc(int size);
import "DPI-C" function void free(chandle ptr); 


