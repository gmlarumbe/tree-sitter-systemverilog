// Section 54.4: Inside

a inside {[0:5], [8:15]};


