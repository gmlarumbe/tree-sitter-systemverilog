// Section 99.2: Struct

struct packed signed {
  int A;
  byte B;
  byte C;
} PackedStruct;               // Signed, 2-state


