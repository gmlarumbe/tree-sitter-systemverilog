module a ();

always @(posedge clk or negedge rst_n) begin end

endmodule
