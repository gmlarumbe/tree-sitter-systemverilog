function void foo();
    this.a.b.c;
endfunction
