module mod ();

  modA #(42) instA (
    .clk (clk),
    .inp(inp )
  );

endmodule
