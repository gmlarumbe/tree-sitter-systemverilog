module mod ();
  wire [W-1:0] a;
endmodule
