packet = packet_in::type_id::create("packet", this);
