module mod ();

  modA instA (
    .clk (clk),
    .inp(inp )
  );

endmodule
