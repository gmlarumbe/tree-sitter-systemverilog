module mod #(
  parameter A=5,
            B=10
)();

endmodule
