`timescale 1ns/ 100ps
