function f;
    left.member = right.member;
endfunction
