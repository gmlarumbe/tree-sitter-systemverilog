module mod;

initial
  if (cond)
    a = 0;
  else if (cond2)
    a = 1;
  else
    a = 2;


endmodule
