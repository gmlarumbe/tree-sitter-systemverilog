module mod ();
  assign z = a | b ^ c & |d == e;
endmodule
