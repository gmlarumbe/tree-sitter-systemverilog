initial begin
    a = foo[b.c.d()];
end

