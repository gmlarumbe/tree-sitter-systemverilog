// Section 55.4: Instantiation

module foo;
//The following is an and-nor, showing an expression in port connection list
nor (F, A&&B, C);        // Not recommended
endmodule

