function void foo();
    super.new();
endfunction
