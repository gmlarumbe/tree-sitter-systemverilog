initial begin
    a.a = b[i][A+B-1:0];
end

