module mod ();
  always_comb foo = bar.baz.bat;
endmodule
