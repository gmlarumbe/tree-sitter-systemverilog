module mod #(
  parameter P1 = 32,
  parameter P2 = P1,
  parameter P3 = (1 * P1)
)();

endmodule
