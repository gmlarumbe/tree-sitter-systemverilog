// Section 20.1: Const

const int A = 1;

class MyClass;
  const int G = 1; // Global constant
  const int I;     // Instance constant
  function new(int x);
    I = 10;        // Instance constant assigned in constructor.
    /*...*/     
  endfunction
endclass


