library rtlLib *.v; // matches all files in the current directory with a .v suffix
library gateLib ./\*.vg; // matches all files in the current directory with a .vg suffix
