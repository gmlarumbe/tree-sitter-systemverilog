// Section 17.1: Comment

// This is a comment
/*
   So is this - across three lines
*/
module ALU /* 8-bit ALU */ (A, B, Opcode, F);
endmodule


