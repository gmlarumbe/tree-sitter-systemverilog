module mod;

initial
  if (cond)
    a = 0;
  else
    a = 1;


endmodule
