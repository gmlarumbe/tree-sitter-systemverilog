assign mst_reqs_o[i].aw = slv_aw_chan.aw;
