function void foo();
    this.fun();
endfunction
