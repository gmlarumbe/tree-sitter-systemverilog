class asdf;

    static function void turn_on_tracing();
        a = init;
        a = init();

        if (!ready)
           a = init();

        tracing = 1;
    endfunction

endclass
