// Section 35.2: Export "DPI-C"

// C:
#include "svdpi.h"
extern void read(int);   // Imported from SystemVerilog


