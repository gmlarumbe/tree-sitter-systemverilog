// Section 18.1: Compilation Unit

bit b;
function void AFunc;
  int b;
  b = $unit::b;     // $unit::b is the one outside
endfunction


