// Section 137.1: Within

property p;
!sig1[*3] within (($fell(sig2)) ##0 !sig2[*5])
endproperty


