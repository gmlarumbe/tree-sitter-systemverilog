function void foo();
    this.super.fun();
endfunction
