function void foo();
    a = init(.arg1(arg1), .arg2(arg2));
endfunction
