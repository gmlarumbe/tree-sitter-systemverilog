// Section 148.1: $unit

initial begin
$unit::semi_global_sig; // Compilation unit name
end

