// Section 45.2: Function

function [15:0][7:0] AFunc(
  int A,                            // A is input by default
  output [15:0][7:0] B, C[15:0]); 
  /*...*/
endfunction


