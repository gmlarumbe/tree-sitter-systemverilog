module a ();

always @* begin end

endmodule
