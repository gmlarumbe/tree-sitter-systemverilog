module a ();

always @(posedge clk) begin end

endmodule
