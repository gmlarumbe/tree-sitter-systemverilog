function f;
    left[i+10] = right[i+10];
endfunction
