// Section 62.2: Library
  
// References any .v source in a project hierarchy, regardless of the directory
// names or structure within it.
// (uncomment the following to use)
// library ProjectLib /usr/design/project//*...*//*.v ;


