`define D(x, y) initial $display("start", x, y)
