initial begin
    a = class1::class2::member1.member2;
end
