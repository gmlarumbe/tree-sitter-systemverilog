function f;
    a = b[1][1];
endfunction
