module test;
    initial begin
        $finish;
    end
endmodule
