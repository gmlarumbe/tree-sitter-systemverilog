`line 10 "bar" 2
