// Section 55.2: Instantiation

//Module instance
Counter U123 (.Clock(Clk), .Reset(Rst), .Count(Q));


