// Section 106.4: Typedef

typedef mailbox #(int) MailBox; // Parameterised mailbox
MailBox MB = new;


