class foo;
endclass
