function void foo();
    a = obj.method();
endfunction
