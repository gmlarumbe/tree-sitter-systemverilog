module mod ();
  assign a = (b == c) ? (d == e) ? (f == g) ? h : i : j : k;
endmodule
