// Section 8.5: Attribute

// Attribute attached to an interface
(*interface_att = 10*) interface Int1; /*...*/ endinterface


