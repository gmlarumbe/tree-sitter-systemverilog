module mod ();

  assign quz = 16'habc;
  assign bar = 6'o42;
  assign foo = 7'b010_1000;
  assign baz = 12'd987654;

endmodule
