  localparam int unsigned AxiIdWidth    = 32'd10;

