function void foo();
    a = super.new();
endfunction
