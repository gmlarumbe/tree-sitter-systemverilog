// Section 74.4: Operators

// Replication operator (or multiple concatenation)
int a = {4{1'b1}};                  // Equivalent to 4'b1111


