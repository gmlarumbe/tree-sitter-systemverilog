function void foo();
    this.in_use[i].get_start_offset();
endfunction
