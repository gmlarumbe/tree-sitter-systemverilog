// Section 104.1: Timeunit

timeunit 100ns;
timeprecision 10ps;


