module test;
    initial begin
        k = $random;
    end
endmodule
