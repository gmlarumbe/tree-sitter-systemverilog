// Section 111.1: Variable

reg a, b, c;
logic [7:0] mem[1:1024], Byte; // Byte is not a memory array
integer i, j, k;
time now;
real r;
shortint ShInt[7];             // Same as ShInt[0:6]
bit[7:0] B;                    // Same as byte B;
logic signed [31:0] L;         // Same as integer L;
byte C = "A";


