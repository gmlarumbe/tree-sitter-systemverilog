class asdf;

    static function void turn_on_tracing();
        init;
        init();

        if (!ready)
           init();

        tracing = 1;
    endfunction

endclass
