`include <bar>
