// Section 74.3: Operators

// Or and , in sensitivity list
always @(A or B, C, D or E)
    begin
    end
