// Section 40.1: Force

force f = a && b;
/*...*/
release f;


