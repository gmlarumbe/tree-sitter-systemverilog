initial begin
    a.a = b[i][A.a+B.b-1:0];
end
