// Section 8.2: Attribute

// Attribute attached to an operator
A = B + (* mode = "cla" *) C; 


