function f;
    left.member.nested[1] = right.member.nested[1];
endfunction
