// Section 2.2: Always

always_comb
  A = B & C;
always_comb
  A <= #10ns B & C;

  
