module a ();

always @(comb1, comb2, comb3, comb4) begin end

endmodule
