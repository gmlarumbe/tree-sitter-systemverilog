module mod ();
  assign a = b == c ? d : e;
endmodule
