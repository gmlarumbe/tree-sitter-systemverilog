typedef shortint unsigned u_shortint_t;
