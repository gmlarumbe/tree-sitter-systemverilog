module mod;

initial begin
  if (cond) begin
    a = 0;
  end
  else if (cond2) begin
    a = 1;
  end
  else begin
    a = 2;
  end
end

endmodule

