class foo extends base_class #(base_type);
endclass
