module mod ();
  assign a = b[3:1];
endmodule
