module foo;

    logic [3:0]           data1;
    logic [3:0][4:0]      data2;
    logic [3:0][4:0][5:0] data3;

endmodule;
