// Section 3.4: Array

// Multiple unpacked dimensions defined in stages using typedef
typedef B8 Mem[0:3];                 // Array of four B8 elements
Mem Mem8[0:7];                       // Array of 8 Mem elements


