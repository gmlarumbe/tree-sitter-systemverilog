module mod (); endmodule
