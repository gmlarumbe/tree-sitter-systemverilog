module mod ();
  assign a = ~|c;
endmodule
