// Section 101.3: Task

// An automatic task with static variables
task automatic Task();
  int VarA1;            // Automatic by default
  static int VarS;      // Static
  automatic int VarA2;  // Automatic
    // /*...*/
endtask


