function void foo();
    this.a.b.c(.arg1(arg1), .arg2(arg2));
endfunction
