module mod;

initial begin
  if (cond) begin
    a = 0;
  end
end

endmodule
