`some_macro(arg1, arg2)
