module mod;

initial
  if (cond)
    a = 0;


endmodule
