function f;
    left.member[1] = right.member[1];
endfunction
