function void foo();
    a = init(arg1, arg2);
endfunction
