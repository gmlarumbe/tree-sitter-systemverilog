// Section 114.2: Wait

// Wait until the sequence seq1 is successfully completed
wait (seq1.triggered)
  $display("Sequence seq1 has completed");


