module a ();

always @(posedge clk, negedge rst_n, signal) begin end

endmodule
