// Section 74.2: Operators

// Assignment to RegA when an event occurs on A or B
@(A, B) RegA = RegB;


