typedef class my_class;
