function void foo();
    if (this.in_use[i+1].get_start_offset() < cfg.start_offset) begin
        ;
    end
endfunction
