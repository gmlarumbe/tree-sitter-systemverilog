/* multi- line comment */
