function f;
    left[1][1:0] = right[1][1:0];
endfunction
