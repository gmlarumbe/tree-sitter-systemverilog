module m
  import mp::*;
`ifdef EX_V
  import mv::*;
`endif
   (
    input logic                              clk,
    input logic                              nrst
   );

endmodule
