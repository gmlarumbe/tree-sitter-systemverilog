function void foo();
    this.in_use[0].get_start_offset();
endfunction
