function f;
    left.member.nested[1][2] = right.member.nested[1][2];
endfunction
