bind cpu: cpu1 fpu_props fpu_rules_1(a, b, c);
