function void foo();
    a = a.b.c();
endfunction
