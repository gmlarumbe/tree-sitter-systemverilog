initial begin
    a = int'(2.0 * 3.0);
    b = shortint'({8'hFA,8'hCE});
    A = cast_t1'(expr_1) + cast_t2'(expr_2);
end

