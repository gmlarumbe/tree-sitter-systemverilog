module mod;

initial begin
  if (cond) begin
    a = 0;
  end
  else begin
    a = 1;
  end
end

endmodule
