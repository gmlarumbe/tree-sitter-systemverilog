module foo # (
    parameter `FOO(arg)
    )();
endmodule
