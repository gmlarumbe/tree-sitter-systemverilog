// Section 54.4: Inside

initial begin
if (a inside {[0:5], [8:15]})
    ;
end


