module mod #(
  parameter A = 5
)(
  output reg [A - 1 : 0] out1,
  output reg [(A - 1): 0] out2
);

endmodule
