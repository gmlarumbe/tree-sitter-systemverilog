package NetsPkg;
  nettype real realNet;
endpackage : NetsPkg
