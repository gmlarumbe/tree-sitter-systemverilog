interface foo;
endinterface
