class driver #(type T=int) extends uvm_component;
  `uvm_component_param_utils(driver #(T));
   //  ...
endclass
