task class_scope::method(input logic in, output logic out);
    foo = foo2;
endtask : method
