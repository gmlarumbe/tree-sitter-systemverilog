module foo;
    and u1 (Q, A, B);
    and #(2.1, 2.8) u2 (Q, A, B);
    and (pull0, strong1) (Q, A, B);
endmodule
