module a_l ();

always @(a or b or c or d) begin end

endmodule
