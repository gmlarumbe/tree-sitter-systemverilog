function f;
    left[A] = right[A];
endfunction
