module mod #()();
endmodule
