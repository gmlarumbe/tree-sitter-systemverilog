// Section 69.1: Name

module foo;
// Legal names
logic A_99_Z;
logic Reset;
logic _54MHz_Clock$;
logic Module;                 // Not the same as 'module'
logic \$%^&*() ;               // Escaped identifier

endmodule
