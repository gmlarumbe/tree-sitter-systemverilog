// Section 106.2: Typedef

typedef struct {byte Addr; byte Data;} Bus; 
Bus Bus1[0:3];                     // Array of structures 


