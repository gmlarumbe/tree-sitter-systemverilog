// Section 116.1: `begin_keywords

`begin_keywords "1364-2001-noconfig"
module design;         // design is a keyword in Verilog-2001
  reg logic;           // logic is a keyword in SystemVerilog
endmodule
`end_keywords


