module foo # (
    parameter `FOO(arg),
    parameter `FOO2(arg2),
    parameter `FOO3,
              identifier = 0,
              other = 1
    )();
endmodule
