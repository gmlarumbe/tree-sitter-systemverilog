module mod ();
  assign a = (
    b + c)
      | &(b
        & 5 );
endmodule
