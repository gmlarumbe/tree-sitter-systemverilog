module x;
    always begin
        a <= {WIDTH{1'b0}};
    end
endmodule
