module mod ();
  assign a = b[0:Param+1];
endmodule
