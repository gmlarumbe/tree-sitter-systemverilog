module mod #(
  parameter A=5,
            B=10,
  parameter C=15,
  localparam D=10
)();

endmodule
