function void foo();
    init(arg1, arg2);
endfunction
