// Section 54.5: Inside

string I;
I inside {["abc":"def"]}       // I between "abc" and "def"


