module mod ();
  assign a = {b,c , d };
endmodule
