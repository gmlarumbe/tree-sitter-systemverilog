module mod ();
  assign a = b[1+Param:0];
endmodule
