// Section 7.2: Associative Array

// Create an array of string, indexed by integers
string Table [*];
Table = '{0:"Zero", 1:"One", 2:"Two", default:"None"};
$display("%s %s", Table[0], Table[3]); // Displays "Zero None"


