initial begin
    class1::class2::member1.member2 = 10;
end
