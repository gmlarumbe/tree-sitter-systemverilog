module mod ();
  assign a = 5;
endmodule
