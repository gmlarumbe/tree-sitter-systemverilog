// Section 78.1: Port

module (A, B, C, D);
  input A;
  inout [7:0] B;
  output [3:0] C, D;
endmodule


