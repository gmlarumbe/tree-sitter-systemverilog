module mod ();
  always_comb foo = bar.baz;
endmodule
