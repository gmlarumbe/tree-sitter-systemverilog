module mod ();

  modA #(.WIDTH(8), .DEPTH(4)) instA (
    .clk (clk)
  );

endmodule
