`default_nettype wire
