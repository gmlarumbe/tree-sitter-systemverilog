function void foo();
    if (a = callbacks.size()) begin
        return;
    end
endfunction
