module foo;
  block u_block (if1.signal, if2.signal);
endmodule : foo
