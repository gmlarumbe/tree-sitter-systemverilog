class foo;
    rand int a = 0;
    randc int b = 1;
endclass
