module mod #(
  parameter type T = logic,
                 Q = bit
)();

endmodule
