// Section 107.1: Union

typedef union packed {
  bit [15:0] i;
  shortint   j;
} Un; 

Un N;
N.j = 0;
	

