// Section 30.1: Do-While

int N = 10;
do
  begin
    /*...*/
    N++;
  end
while (N < 100);


