function void foo();
    if (this.in_use[0].get_start_offset() < cfg.start_offset) begin
        ;
    end
endfunction
