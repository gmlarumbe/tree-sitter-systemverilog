include rtlLib *.v;
include gateLib ./\*.vg;
