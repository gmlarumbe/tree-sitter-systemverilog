module foo;
    specify
        specparam PATHPULSE$ = (0.5);
    endspecify
endmodule
