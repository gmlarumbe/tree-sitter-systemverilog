// Section 144.1: $root

initial begin
$root.MyModule.U1; // Absolute name
end

