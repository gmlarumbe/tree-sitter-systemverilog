module mod ();

  modA instA (clk, inp);

endmodule
