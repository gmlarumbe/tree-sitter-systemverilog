function void foo();
    obj.method();
endfunction
