function void foo();
    a = this.a.b.c;
endfunction
