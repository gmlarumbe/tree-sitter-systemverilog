function void foo();
    a.b.c();
endfunction
