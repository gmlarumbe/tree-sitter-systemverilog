module test;
    initial begin
        $print("%d, %d, %d", a, b, c);
    end
endmodule
