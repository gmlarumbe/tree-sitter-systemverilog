// Section 3.3: Array

// Multiple packed dimensions defined in stages using typedef
typedef bit [0:7] B8;
B8 [0:15] B8_16;                     // [0:7] varies most rapidly


