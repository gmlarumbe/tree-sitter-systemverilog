module x;
    always begin
        a <= {{1'b0,1'b0}};
    end
endmodule
