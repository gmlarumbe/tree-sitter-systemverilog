// Section 8.4: Attribute

// Attribute attached to a conditional operator 
A = B ? (* no_glitch *) C : D; 


