function void foo();
    if(!this.randomize()) begin
        return;
    end
endfunction
