function void foo();
    if (this.in_use[i].get_start_offset() < cfg.start_offset) begin
        ;
    end
endfunction
