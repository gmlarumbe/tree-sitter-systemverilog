// Section 78.2: Port

module FF8(
  input Clk, Reset,
  input reg [7:0] D,
  output reg [7:0] Q = 8'b0); // Declare and initialize reg
endmodule

