module foo;
    my_and u1 (Q, A, B);
    my_and #(2.1, 2.8) u2 (Q, A, B);
    my_and (Q, A, B);
    my_and (pull0, strong1) (Q, A, B);
endmodule
