module mod ();

  modA instA ();

endmodule
