// Section 6.1: Assign

//Continuous assignment
wire cout, cin;
wire [31:0] sum, a, b;

assign {cout, sum} = a + b + cin;


