bind cr_unit range r1(c_clk,c_en,v_low,(in1&&in2));
