initial begin
  string a = """
  a, b, c, "xy"
  """;
end
