initial begin
    string inst_name;
    inst_name = {slash_or_blank,
                 cntxt.get_full_name(),
                 separator,
                 inst_name,
                 close_or_blank};
end


