module abc ();

always_comb
if (a) begin
  a = b;
end

endmodule
