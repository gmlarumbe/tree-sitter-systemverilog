function f;
    left.member.nested[1][2][1:0] = right.member.nested[1][2][1:0];
endfunction
