class foo;
    function new ();
    endfunction : new
endclass
