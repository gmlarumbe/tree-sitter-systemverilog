function void foo;
    a = class_type::method();
endfunction
