// Section 3.2: Array

// Reading and writing a variable slice of the array
A[x+:c] = B[y+:c];                   // c must be constant


