// Section 133.1: Property

property P;
  (a ##1 b) |-> (d ##1 e);
endproperty


