initial begin
    mem_n[8'(trans_id_i[i])-1].sbe.valid = 1'b1;
end
