// Section 106.1: Typedef

typedef enum {True, False} Bool;
Bool Var; 


