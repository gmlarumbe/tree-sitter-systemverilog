function f;
    a = b[1];
endfunction
