// Section 139.1: $display and $write

$display("Illegal opcode %h in %m at %t",
          Opcode, $realtime);

$writeh("Variable values (hex.): ",
          reg1,, reg2,, reg3,, reg4,"\n");


