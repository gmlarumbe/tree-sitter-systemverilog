// Section 76.3: Parameter

// Typed parameters
parameter integer Size = 1;


