typedef enum int {RED, YELLOW, BLUE} light_e;
typedef struct {
    logic  element_1;
    logic  element_2;
    } my_struct_t;
