function void foo();
    if(a = !this.randomize()) begin
        return;
    end
endfunction
