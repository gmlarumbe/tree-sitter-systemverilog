class foo;

    function void foo;
    endfunction

    task foo;
    endtask

endclass
