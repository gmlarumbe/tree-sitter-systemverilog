function foo;
   class_id.attribute = value;
endfunction
