class foo #(int N=1, int P=2);
endclass
