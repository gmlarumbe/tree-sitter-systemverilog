module mod ();
  assign a = b & c;
endmodule
