// Section 76.5: Parameter

// Parameter dependence
parameter WordSize = 16, MemSize = WordSize*1024;


