function void foo;
  `MY_MACRO.identifier[0].member = 0;
endfunction
