function f;
    left[A][1:0] = right[A][1:0];
endfunction
